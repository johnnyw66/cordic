
module  circle256_2_28  (
	input clk,
	input  [7:0] cangle,
	output reg [WIDTH-1:0] rangle
);

parameter WIDTH = 32 ;


// Fixed point radian Angles (2:28)
//   (index * 2.0 * math.pi / 256) * (1 << 32)

always @(posedge clk)
begin
  case(cangle)
      8'd00 : rangle <= 32'b0000000000000000000000000000000 ;
      8'd01 : rangle <= 32'b0000000011001001000011111101101 ;
      8'd02 : rangle <= 32'b0000000110010010000111111011010 ;
      8'd03 : rangle <= 32'b0000001001011011001011111000111 ;
      8'd04 : rangle <= 32'b0000001100100100001111110110101 ;
      8'd05 : rangle <= 32'b0000001111101101010011110100010 ;
      8'd06 : rangle <= 32'b0000010010110110010111110001111 ;
      8'd07 : rangle <= 32'b0000010101111111011011101111101 ;
      8'd08 : rangle <= 32'b0000011001001000011111101101010 ;
      8'd09 : rangle <= 32'b0000011100010001100011101010111 ;
      8'd10 : rangle <= 32'b0000011111011010100111101000101 ;
      8'd11 : rangle <= 32'b0000100010100011101011100110010 ;
      8'd12 : rangle <= 32'b0000100101101100101111100011111 ;
      8'd13 : rangle <= 32'b0000101000110101110011100001101 ;
      8'd14 : rangle <= 32'b0000101011111110110111011111010 ;
      8'd15 : rangle <= 32'b0000101111000111111011011100111 ;
      8'd16 : rangle <= 32'b0000110010010000111111011010101 ;
      8'd17 : rangle <= 32'b0000110101011010000011011000010 ;
      8'd18 : rangle <= 32'b0000111000100011000111010101111 ;
      8'd19 : rangle <= 32'b0000111011101100001011010011101 ;
      8'd20 : rangle <= 32'b0000111110110101001111010001010 ;
      8'd21 : rangle <= 32'b0001000001111110010011001110111 ;
      8'd22 : rangle <= 32'b0001000101000111010111001100100 ;
      8'd23 : rangle <= 32'b0001001000010000011011001010010 ;
      8'd24 : rangle <= 32'b0001001011011001011111000111111 ;
      8'd25 : rangle <= 32'b0001001110100010100011000101100 ;
      8'd26 : rangle <= 32'b0001010001101011100111000011010 ;
      8'd27 : rangle <= 32'b0001010100110100101011000000111 ;
      8'd28 : rangle <= 32'b0001010111111101101110111110100 ;
      8'd29 : rangle <= 32'b0001011011000110110010111100010 ;
      8'd30 : rangle <= 32'b0001011110001111110110111001111 ;
      8'd31 : rangle <= 32'b0001100001011000111010110111100 ;
      8'd32 : rangle <= 32'b0001100100100001111110110101010 ;
      8'd33 : rangle <= 32'b0001100111101011000010110010111 ;
      8'd34 : rangle <= 32'b0001101010110100000110110000100 ;
      8'd35 : rangle <= 32'b0001101101111101001010101110010 ;
      8'd36 : rangle <= 32'b0001110001000110001110101011111 ;
      8'd37 : rangle <= 32'b0001110100001111010010101001100 ;
      8'd38 : rangle <= 32'b0001110111011000010110100111010 ;
      8'd39 : rangle <= 32'b0001111010100001011010100100111 ;
      8'd40 : rangle <= 32'b0001111101101010011110100010100 ;
      8'd41 : rangle <= 32'b0010000000110011100010100000001 ;
      8'd42 : rangle <= 32'b0010000011111100100110011101111 ;
      8'd43 : rangle <= 32'b0010000111000101101010011011100 ;
      8'd44 : rangle <= 32'b0010001010001110101110011001001 ;
      8'd45 : rangle <= 32'b0010001101010111110010010110111 ;
      8'd46 : rangle <= 32'b0010010000100000110110010100100 ;
      8'd47 : rangle <= 32'b0010010011101001111010010010001 ;
      8'd48 : rangle <= 32'b0010010110110010111110001111111 ;
      8'd49 : rangle <= 32'b0010011001111100000010001101100 ;
      8'd50 : rangle <= 32'b0010011101000101000110001011001 ;
      8'd51 : rangle <= 32'b0010100000001110001010001000111 ;
      8'd52 : rangle <= 32'b0010100011010111001110000110100 ;
      8'd53 : rangle <= 32'b0010100110100000010010000100001 ;
      8'd54 : rangle <= 32'b0010101001101001010110000001111 ;
      8'd55 : rangle <= 32'b0010101100110010011001111111100 ;
      8'd56 : rangle <= 32'b0010101111111011011101111101001 ;
      8'd57 : rangle <= 32'b0010110011000100100001111010111 ;
      8'd58 : rangle <= 32'b0010110110001101100101111000100 ;
      8'd59 : rangle <= 32'b0010111001010110101001110110001 ;
      8'd60 : rangle <= 32'b0010111100011111101101110011110 ;
      8'd61 : rangle <= 32'b0010111111101000110001110001100 ;
      8'd62 : rangle <= 32'b0011000010110001110101101111001 ;
      8'd63 : rangle <= 32'b0011000101111010111001101100110 ;
      8'd64 : rangle <= 32'b0011001001000011111101101010100 ;
      8'd65 : rangle <= 32'b0011001100001101000001101000001 ;
      8'd66 : rangle <= 32'b0011001111010110000101100101110 ;
      8'd67 : rangle <= 32'b0011010010011111001001100011100 ;
      8'd68 : rangle <= 32'b0011010101101000001101100001001 ;
      8'd69 : rangle <= 32'b0011011000110001010001011110110 ;
      8'd70 : rangle <= 32'b0011011011111010010101011100100 ;
      8'd71 : rangle <= 32'b0011011111000011011001011010001 ;
      8'd72 : rangle <= 32'b0011100010001100011101010111110 ;
      8'd73 : rangle <= 32'b0011100101010101100001010101100 ;
      8'd74 : rangle <= 32'b0011101000011110100101010011001 ;
      8'd75 : rangle <= 32'b0011101011100111101001010000110 ;
      8'd76 : rangle <= 32'b0011101110110000101101001110100 ;
      8'd77 : rangle <= 32'b0011110001111001110001001100001 ;
      8'd78 : rangle <= 32'b0011110101000010110101001001110 ;
      8'd79 : rangle <= 32'b0011111000001011111001000111100 ;
      8'd80 : rangle <= 32'b0011111011010100111101000101001 ;
      8'd81 : rangle <= 32'b0011111110011110000001000010110 ;
      8'd82 : rangle <= 32'b0100000001100111000101000000011 ;
      8'd83 : rangle <= 32'b0100000100110000001000111110001 ;
      8'd84 : rangle <= 32'b0100000111111001001100111011110 ;
      8'd85 : rangle <= 32'b0100001011000010010000111001011 ;
      8'd86 : rangle <= 32'b0100001110001011010100110111001 ;
      8'd87 : rangle <= 32'b0100010001010100011000110100110 ;
      8'd88 : rangle <= 32'b0100010100011101011100110010011 ;
      8'd89 : rangle <= 32'b0100010111100110100000110000001 ;
      8'd90 : rangle <= 32'b0100011010101111100100101101110 ;
      8'd91 : rangle <= 32'b0100011101111000101000101011011 ;
      8'd92 : rangle <= 32'b0100100001000001101100101001001 ;
      8'd93 : rangle <= 32'b0100100100001010110000100110110 ;
      8'd94 : rangle <= 32'b0100100111010011110100100100011 ;
      8'd95 : rangle <= 32'b0100101010011100111000100010001 ;
      8'd96 : rangle <= 32'b0100101101100101111100011111110 ;
      8'd97 : rangle <= 32'b0100110000101111000000011101011 ;
      8'd98 : rangle <= 32'b0100110011111000000100011011001 ;
      8'd99 : rangle <= 32'b0100110111000001001000011000110 ;
      8'd100 : rangle <= 32'b0100111010001010001100010110011 ;
      8'd101 : rangle <= 32'b0100111101010011010000010100000 ;
      8'd102 : rangle <= 32'b0101000000011100010100010001110 ;
      8'd103 : rangle <= 32'b0101000011100101011000001111011 ;
      8'd104 : rangle <= 32'b0101000110101110011100001101000 ;
      8'd105 : rangle <= 32'b0101001001110111100000001010110 ;
      8'd106 : rangle <= 32'b0101001101000000100100001000011 ;
      8'd107 : rangle <= 32'b0101010000001001101000000110000 ;
      8'd108 : rangle <= 32'b0101010011010010101100000011110 ;
      8'd109 : rangle <= 32'b0101010110011011110000000001011 ;
      8'd110 : rangle <= 32'b0101011001100100110011111111000 ;
      8'd111 : rangle <= 32'b0101011100101101110111111100110 ;
      8'd112 : rangle <= 32'b0101011111110110111011111010011 ;
      8'd113 : rangle <= 32'b0101100010111111111111111000000 ;
      8'd114 : rangle <= 32'b0101100110001001000011110101110 ;
      8'd115 : rangle <= 32'b0101101001010010000111110011011 ;
      8'd116 : rangle <= 32'b0101101100011011001011110001000 ;
      8'd117 : rangle <= 32'b0101101111100100001111101110110 ;
      8'd118 : rangle <= 32'b0101110010101101010011101100011 ;
      8'd119 : rangle <= 32'b0101110101110110010111101010000 ;
      8'd120 : rangle <= 32'b0101111000111111011011100111101 ;
      8'd121 : rangle <= 32'b0101111100001000011111100101011 ;
      8'd122 : rangle <= 32'b0101111111010001100011100011000 ;
      8'd123 : rangle <= 32'b0110000010011010100111100000101 ;
      8'd124 : rangle <= 32'b0110000101100011101011011110011 ;
      8'd125 : rangle <= 32'b0110001000101100101111011100000 ;
      8'd126 : rangle <= 32'b0110001011110101110011011001101 ;
      8'd127 : rangle <= 32'b0110001110111110110111010111011 ;
      8'd128 : rangle <= 32'b0110010010000111111011010101000 ;
      8'd129 : rangle <= 32'b0110010101010000111111010010101 ;
      8'd130 : rangle <= 32'b0110011000011010000011010000011 ;
      8'd131 : rangle <= 32'b0110011011100011000111001110000 ;
      8'd132 : rangle <= 32'b0110011110101100001011001011101 ;
      8'd133 : rangle <= 32'b0110100001110101001111001001011 ;
      8'd134 : rangle <= 32'b0110100100111110010011000111000 ;
      8'd135 : rangle <= 32'b0110101000000111010111000100101 ;
      8'd136 : rangle <= 32'b0110101011010000011011000010011 ;
      8'd137 : rangle <= 32'b0110101110011001011111000000000 ;
      8'd138 : rangle <= 32'b0110110001100010100010111101101 ;
      8'd139 : rangle <= 32'b0110110100101011100110111011011 ;
      8'd140 : rangle <= 32'b0110110111110100101010111001000 ;
      8'd141 : rangle <= 32'b0110111010111101101110110110101 ;
      8'd142 : rangle <= 32'b0110111110000110110010110100010 ;
      8'd143 : rangle <= 32'b0111000001001111110110110010000 ;
      8'd144 : rangle <= 32'b0111000100011000111010101111101 ;
      8'd145 : rangle <= 32'b0111000111100001111110101101010 ;
      8'd146 : rangle <= 32'b0111001010101011000010101011000 ;
      8'd147 : rangle <= 32'b0111001101110100000110101000101 ;
      8'd148 : rangle <= 32'b0111010000111101001010100110010 ;
      8'd149 : rangle <= 32'b0111010100000110001110100100000 ;
      8'd150 : rangle <= 32'b0111010111001111010010100001101 ;
      8'd151 : rangle <= 32'b0111011010011000010110011111010 ;
      8'd152 : rangle <= 32'b0111011101100001011010011101000 ;
      8'd153 : rangle <= 32'b0111100000101010011110011010101 ;
      8'd154 : rangle <= 32'b0111100011110011100010011000010 ;
      8'd155 : rangle <= 32'b0111100110111100100110010110000 ;
      8'd156 : rangle <= 32'b0111101010000101101010010011101 ;
      8'd157 : rangle <= 32'b0111101101001110101110010001010 ;
      8'd158 : rangle <= 32'b0111110000010111110010001111000 ;
      8'd159 : rangle <= 32'b0111110011100000110110001100101 ;
      8'd160 : rangle <= 32'b0111110110101001111010001010010 ;
      8'd161 : rangle <= 32'b0111111001110010111110000111111 ;
      8'd162 : rangle <= 32'b0111111100111100000010000101101 ;
      8'd163 : rangle <= 32'b1000000000000101000110000011010 ;
      8'd164 : rangle <= 32'b1000000011001110001010000000111 ;
      8'd165 : rangle <= 32'b1000000110010111001101111110101 ;
      8'd166 : rangle <= 32'b1000001001100000010001111100010 ;
      8'd167 : rangle <= 32'b1000001100101001010101111001111 ;
      8'd168 : rangle <= 32'b1000001111110010011001110111101 ;
      8'd169 : rangle <= 32'b1000010010111011011101110101010 ;
      8'd170 : rangle <= 32'b1000010110000100100001110010111 ;
      8'd171 : rangle <= 32'b1000011001001101100101110000101 ;
      8'd172 : rangle <= 32'b1000011100010110101001101110010 ;
      8'd173 : rangle <= 32'b1000011111011111101101101011111 ;
      8'd174 : rangle <= 32'b1000100010101000110001101001101 ;
      8'd175 : rangle <= 32'b1000100101110001110101100111010 ;
      8'd176 : rangle <= 32'b1000101000111010111001100100111 ;
      8'd177 : rangle <= 32'b1000101100000011111101100010101 ;
      8'd178 : rangle <= 32'b1000101111001101000001100000010 ;
      8'd179 : rangle <= 32'b1000110010010110000101011101111 ;
      8'd180 : rangle <= 32'b1000110101011111001001011011100 ;
      8'd181 : rangle <= 32'b1000111000101000001101011001010 ;
      8'd182 : rangle <= 32'b1000111011110001010001010110111 ;
      8'd183 : rangle <= 32'b1000111110111010010101010100100 ;
      8'd184 : rangle <= 32'b1001000010000011011001010010010 ;
      8'd185 : rangle <= 32'b1001000101001100011101001111111 ;
      8'd186 : rangle <= 32'b1001001000010101100001001101100 ;
      8'd187 : rangle <= 32'b1001001011011110100101001011010 ;
      8'd188 : rangle <= 32'b1001001110100111101001001000111 ;
      8'd189 : rangle <= 32'b1001010001110000101101000110100 ;
      8'd190 : rangle <= 32'b1001010100111001110001000100010 ;
      8'd191 : rangle <= 32'b1001011000000010110101000001111 ;
      8'd192 : rangle <= 32'b1001011011001011111000111111100 ;
      8'd193 : rangle <= 32'b1001011110010100111100111101010 ;
      8'd194 : rangle <= 32'b1001100001011110000000111010111 ;
      8'd195 : rangle <= 32'b1001100100100111000100111000100 ;
      8'd196 : rangle <= 32'b1001100111110000001000110110010 ;
      8'd197 : rangle <= 32'b1001101010111001001100110011111 ;
      8'd198 : rangle <= 32'b1001101110000010010000110001100 ;
      8'd199 : rangle <= 32'b1001110001001011010100101111010 ;
      8'd200 : rangle <= 32'b1001110100010100011000101100111 ;
      8'd201 : rangle <= 32'b1001110111011101011100101010100 ;
      8'd202 : rangle <= 32'b1001111010100110100000101000001 ;
      8'd203 : rangle <= 32'b1001111101101111100100100101111 ;
      8'd204 : rangle <= 32'b1010000000111000101000100011100 ;
      8'd205 : rangle <= 32'b1010000100000001101100100001001 ;
      8'd206 : rangle <= 32'b1010000111001010110000011110111 ;
      8'd207 : rangle <= 32'b1010001010010011110100011100100 ;
      8'd208 : rangle <= 32'b1010001101011100111000011010001 ;
      8'd209 : rangle <= 32'b1010010000100101111100010111111 ;
      8'd210 : rangle <= 32'b1010010011101111000000010101100 ;
      8'd211 : rangle <= 32'b1010010110111000000100010011001 ;
      8'd212 : rangle <= 32'b1010011010000001001000010000111 ;
      8'd213 : rangle <= 32'b1010011101001010001100001110100 ;
      8'd214 : rangle <= 32'b1010100000010011010000001100001 ;
      8'd215 : rangle <= 32'b1010100011011100010100001001111 ;
      8'd216 : rangle <= 32'b1010100110100101011000000111100 ;
      8'd217 : rangle <= 32'b1010101001101110011100000101001 ;
      8'd218 : rangle <= 32'b1010101100110111100000000010111 ;
      8'd219 : rangle <= 32'b1010110000000000100100000000100 ;
      8'd220 : rangle <= 32'b1010110011001001100111111110001 ;
      8'd221 : rangle <= 32'b1010110110010010101011111011110 ;
      8'd222 : rangle <= 32'b1010111001011011101111111001100 ;
      8'd223 : rangle <= 32'b1010111100100100110011110111001 ;
      8'd224 : rangle <= 32'b1010111111101101110111110100110 ;
      8'd225 : rangle <= 32'b1011000010110110111011110010100 ;
      8'd226 : rangle <= 32'b1011000101111111111111110000001 ;
      8'd227 : rangle <= 32'b1011001001001001000011101101110 ;
      8'd228 : rangle <= 32'b1011001100010010000111101011100 ;
      8'd229 : rangle <= 32'b1011001111011011001011101001001 ;
      8'd230 : rangle <= 32'b1011010010100100001111100110110 ;
      8'd231 : rangle <= 32'b1011010101101101010011100100100 ;
      8'd232 : rangle <= 32'b1011011000110110010111100010001 ;
      8'd233 : rangle <= 32'b1011011011111111011011011111110 ;
      8'd234 : rangle <= 32'b1011011111001000011111011101100 ;
      8'd235 : rangle <= 32'b1011100010010001100011011011001 ;
      8'd236 : rangle <= 32'b1011100101011010100111011000110 ;
      8'd237 : rangle <= 32'b1011101000100011101011010110100 ;
      8'd238 : rangle <= 32'b1011101011101100101111010100001 ;
      8'd239 : rangle <= 32'b1011101110110101110011010001110 ;
      8'd240 : rangle <= 32'b1011110001111110110111001111011 ;
      8'd241 : rangle <= 32'b1011110101000111111011001101001 ;
      8'd242 : rangle <= 32'b1011111000010000111111001010110 ;
      8'd243 : rangle <= 32'b1011111011011010000011001000011 ;
      8'd244 : rangle <= 32'b1011111110100011000111000110001 ;
      8'd245 : rangle <= 32'b1100000001101100001011000011110 ;
      8'd246 : rangle <= 32'b1100000100110101001111000001011 ;
      8'd247 : rangle <= 32'b1100000111111110010010111111001 ;
      8'd248 : rangle <= 32'b1100001011000111010110111100110 ;
      8'd249 : rangle <= 32'b1100001110010000011010111010011 ;
      8'd250 : rangle <= 32'b1100010001011001011110111000001 ;
      8'd251 : rangle <= 32'b1100010100100010100010110101110 ;
      8'd252 : rangle <= 32'b1100010111101011100110110011011 ;
      8'd253 : rangle <= 32'b1100011010110100101010110001001 ;
      8'd254 : rangle <= 32'b1100011101111101101110101110110 ;
      8'd255 : rangle <= 32'b1100100001000110110010101100011 ;
  endcase
end

endmodule
